��
l��F� j�P.�M�.�}q (X   protocol_versionqM�X   little_endianq�X
   type_sizesq}q(X   shortqKX   intqKX   longqKuu.�ccollections
OrderedDict
q )Rq(X   weightqctorch._utils
_rebuild_tensor_v2
q((X   storageqctorch
FloatStorage
qX   93942839980096qX   cpuqKNtqQK KK�q	KK�q
�h )RqtqRqX   biasqh((hhX   93942840064016qhKNtqQK K�qK�q�h )RqtqRqu}qX	   _metadataqh )RqX    q}qX   versionqKsssb.�]q (X   93942839980096qX   93942840064016qe.       �z��gr�@�������       `�